module tb_top;

	reg [3:0] a, b;
	wire [3:0] sum;
	wire [7:0] product;

  top_dut dut1 (.a(a), .b(b), .sum(sum), .product(product)); 

	initial begin

	$dumpfile("dump.vcd");
	$dumpvars(0, tb_top);

        // Mensajes de seguimiento
    $display("Tiempo | a b | sum product");
    $monitor("%4t | %d %d | %d %d", 
              $time, tb_top.a, tb_top.b, tb_top.sum, tb_top.product);
 
		#50 $finish;
 
	end
endmodule
